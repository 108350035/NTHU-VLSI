************************************************************************
* auCdl Netlist:
* 
* Library Name:  mylib
* Top Cell Name: NAND2
* View Name:     schematic
* Netlisted on:  Feb 17 10:39:22 2025
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: mylib
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Vout
*.PININFO A:I B:I VDD:I VSS:I Vout:O
MM1 Vout A VDD VDD p_18 W=1u L=180n
MM0 Vout B VDD VDD p_18 W=1u L=180n
MM3 net15 B VSS VSS n_18 W=0.5u L=180n
MM2 Vout A net15 VSS n_18 W=0.5u L=180n
.ENDS

