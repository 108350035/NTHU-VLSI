************************************************************************
* auCdl Netlist:
* 
* Library Name:  mylib
* Top Cell Name: IV_curves_N
* View Name:     schematic
* Netlisted on:  Feb 15 21:23:19 2025
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: mylib
* Cell Name:    IV_curves_N
* View Name:    schematic
************************************************************************

.SUBCKT IV_curves_N Vds Vgs Vss
*.PININFO Vds:I Vgs:I Vss:I
MM0 Vds Vgs Vss Vss n_18 W=500.0n L=180.00n m=1
.ENDS

