* File: /home/IC/lab6/BUF/buf.pex.spi
* Created: Sat Feb 22 21:29:41 2025
* Program "Calibre xRC"
* Version "v2019.3_15.11"
* 
.include "/home/IC/lab6/BUF/buf.pex.spi.pex"
.subckt BUF  A OUT VSS VDD
* 
* VDD	VDD
* VSS	VSS
* OUT	OUT
* A	A
mXI3.MM1 N_NET07_XI3.MM1_d N_A_XI3.MM1_g N_VSS_XI3.MM1_s N_VSS_XI3.MM1_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.5e-13 PD=1.48e-06 PS=1.5e-06
MM0 N_OUT_MM0_d N_NET07_MM0_g N_VSS_MM0_s N_VSS_XI3.MM1_b N_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXI3.MM0 N_NET07_XI3.MM0_d N_A_XI3.MM0_g N_VDD_XI3.MM0_s N_VDD_XI3.MM0_b P_18
+ L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
MM1 N_OUT_MM1_d N_NET07_MM1_g N_VDD_MM1_s N_VDD_XI3.MM0_b P_18 L=1.8e-07
+ W=2.67e-06 AD=1.3083e-12 AS=1.3083e-12 PD=3.65e-06 PS=3.65e-06
*
.include "/home/IC/lab6/BUF/buf.pex.spi.BUF.pxi"
*
.ends
*
*
