* File: /home/IC/lab6/NAND2/nand2.pex.spi
* Created: Sun Feb 23 11:15:29 2025
* Program "Calibre xRC"
* Version "v2019.3_15.11"
* 
.include "/home/IC/lab6/NAND2/nand2.pex.spi.pex"
.subckt NAND2  A VOUT B VSS VDD
* 
* VDD	VDD
* VSS	VSS
* B	B
* VOUT	VOUT
* A	A
MM2 N_NET15_MM2_d N_A_MM2_g N_VSS_MM2_s N_VSS_MM2_b N_18 L=1.8e-07 W=2e-06
+ AD=5.1e-13 AS=9.8e-13 PD=5.1e-07 PS=2.98e-06
MM3 N_VOUT_MM3_d N_B_MM3_g N_NET15_MM3_s N_VSS_MM2_b N_18 L=1.8e-07 W=2e-06
+ AD=1.02e-12 AS=5.1e-13 PD=3.02e-06 PS=5.1e-07
MM1 N_VOUT_MM1_d N_A_MM1_g N_VDD_MM1_s N_VDD_MM1_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
MM0 N_VOUT_MM0_d N_B_MM0_g N_VDD_MM0_s N_VDD_MM1_b P_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=5.1e-13 PD=5.1e-07 PS=2.02e-06
*
.include "/home/IC/lab6/NAND2/nand2.pex.spi.NAND2.pxi"
*
.ends
*
*
