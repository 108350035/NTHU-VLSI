* File: /home/IC/lab6/BCLKGEN/bclkgen.pex.spi
* Created: Mon Feb 24 09:57:49 2025
* Program "Calibre xRC"
* Version "v2019.3_15.11"
* 
.include "/home/IC/lab6/BCLKGEN/bclkgen.pex.spi.pex"
.subckt Bclkgen  TRIGGER CLKOUT VSS VDD
* 
* VDD	VDD
* VSS	VSS
* CLKOUT	CLKOUT
* TRIGGER	TRIGGER
mXI0.MM2 N_XI0.NET15_XI0.MM2_d N_TRIGGER_XI0.MM2_g N_VSS_XI0.MM2_s
+ N_VSS_XI3.MM1_b N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=9.8e-13 PD=5.1e-07
+ PS=2.98e-06
mXI0.MM3 N_NET16_XI0.MM3_d N_NET10_XI0.MM3_g N_XI0.NET15_XI0.MM3_s
+ N_VSS_XI3.MM1_b N_18 L=1.8e-07 W=2e-06 AD=1.02e-12 AS=5.1e-13 PD=3.02e-06
+ PS=5.1e-07
mXI7.MM4 N_XI7.NET07_XI7.MM4_d N_NET10_XI7.MM4_g N_VSS_XI7.MM4_s N_VSS_XI3.MM1_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.5e-13 PD=1.48e-06 PS=1.5e-06
mXI7.MM0 N_CLKOUT_XI7.MM0_d N_XI7.NET07_XI7.MM0_g N_VSS_XI7.MM0_s
+ N_VSS_XI3.MM1_b N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06
+ PS=1.98e-06
mXI0.MM1 N_NET16_XI0.MM1_d N_TRIGGER_XI0.MM1_g N_VDD_XI0.MM1_s N_VDD_XI3.MM0_b
+ P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI0.MM0 N_NET16_XI0.MM0_d N_NET10_XI0.MM0_g N_VDD_XI0.MM0_s N_VDD_XI3.MM0_b
+ P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=5.1e-13 PD=5.1e-07 PS=2.02e-06
mXI7.MM5 N_XI7.NET07_XI7.MM5_d N_NET10_XI7.MM5_g N_VDD_XI7.MM5_s N_VDD_XI3.MM0_b
+ P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXI7.MM1 N_CLKOUT_XI7.MM1_d N_XI7.NET07_XI7.MM1_g N_VDD_XI7.MM1_s
+ N_VDD_XI3.MM0_b P_18 L=1.8e-07 W=2.67e-06 AD=1.3083e-12 AS=1.3083e-12
+ PD=3.65e-06 PS=3.65e-06
mXI3.MM1 N_NET21_XI3.MM1_d N_NET16_XI3.MM1_g N_VSS_XI3.MM1_s N_VSS_XI3.MM1_b
+ N_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI3.MM0 N_NET21_XI3.MM0_d N_NET16_XI3.MM0_g N_VDD_XI3.MM0_s N_VDD_XI3.MM0_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06
mXI2.MM1 N_NET15_XI2.MM1_d N_NET21_XI2.MM1_g N_VSS_XI2.MM1_s N_VSS_XI3.MM1_b
+ N_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI2.MM0 N_NET15_XI2.MM0_d N_NET21_XI2.MM0_g N_VDD_XI2.MM0_s N_VDD_XI3.MM0_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06
mXI4.MM1 N_NET14_XI4.MM1_d N_NET15_XI4.MM1_g N_VSS_XI4.MM1_s N_VSS_XI3.MM1_b
+ N_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI4.MM0 N_NET14_XI4.MM0_d N_NET15_XI4.MM0_g N_VDD_XI4.MM0_s N_VDD_XI3.MM0_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06
mXI5.MM1 N_NET13_XI5.MM1_d N_NET14_XI5.MM1_g N_VSS_XI5.MM1_s N_VSS_XI3.MM1_b
+ N_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI5.MM0 N_NET13_XI5.MM0_d N_NET14_XI5.MM0_g N_VDD_XI5.MM0_s N_VDD_XI3.MM0_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06
mXI6.MM1 N_NET12_XI6.MM1_d N_NET13_XI6.MM1_g N_VSS_XI6.MM1_s N_VSS_XI3.MM1_b
+ N_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI6.MM0 N_NET12_XI6.MM0_d N_NET13_XI6.MM0_g N_VDD_XI6.MM0_s N_VDD_XI3.MM0_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06
mXI1.MM1 N_NET10_XI1.MM1_d N_NET12_XI1.MM1_g N_VSS_XI1.MM1_s N_VSS_XI3.MM1_b
+ N_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI1.MM0 N_NET10_XI1.MM0_d N_NET12_XI1.MM0_g N_VDD_XI1.MM0_s N_VDD_XI3.MM0_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06
*
.include "/home/IC/lab6/BCLKGEN/bclkgen.pex.spi.BCLKGEN.pxi"
*
.ends
*
*
