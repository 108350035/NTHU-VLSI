* File: /home/IC/lab6/INV/inv.pex.spi
* Created: Sun Feb 23 20:10:10 2025
* Program "Calibre xRC"
* Version "v2019.3_15.11"
* 
.include "/home/IC/lab6/INV/inv.pex.spi.pex"
.subckt INV  A OUT VSS VDD
* 
* VDD	VDD
* VSS	VSS
* OUT	OUT
* A	A
MM1 N_OUT_MM1_d N_A_MM1_g N_VSS_MM1_s N_VSS_MM1_b N_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
MM0 N_OUT_MM0_d N_A_MM0_g N_VDD_MM0_s N_VDD_MM0_b P_18 L=1.8e-07 W=3e-06
+ AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06
*
.include "/home/IC/lab6/INV/inv.pex.spi.INV.pxi"
*
.ends
*
*
