************************************************************************
* auCdl Netlist:
* 
* Library Name:  mylib
* Top Cell Name: INV
* View Name:     schematic
* Netlisted on:  Feb 15 15:20:17 2025
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: mylib
* Cell Name:    INV
* View Name:    schematic
************************************************************************

.SUBCKT INV A Out VDD VSS
*.PININFO A:I Out:O VDD:I VSS:I
MM1 Out A VSS VSS n_18 W=1u L=180.00n
MM0 Out A VDD VDD p_18 W=2u L=180.00n
.ENDS

