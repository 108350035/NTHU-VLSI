* File: /home/IC/lab6/CLKGEN/clkgen.pex.spi
* Created: Sun Feb 23 20:24:08 2025
* Program "Calibre xRC"
* Version "v2019.3_15.11"
* 
.include "/home/IC/lab6/CLKGEN/clkgen.pex.spi.pex"
.subckt clkgen  A CLKOUT VSS VDD
* 
* VDD	VDD
* VSS	VSS
* CLKOUT	CLKOUT
* A	A
mXI18.MM2 N_XI18.NET15_XI18.MM2_d N_A_XI18.MM2_g N_VSS_XI18.MM2_s
+ N_VSS_XI20.MM1_b N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=9.8e-13 PD=5.1e-07
+ PS=2.98e-06
mXI18.MM3 N_NET27_XI18.MM3_d N_CLKOUT_XI18.MM3_g N_XI18.NET15_XI18.MM3_s
+ N_VSS_XI20.MM1_b N_18 L=1.8e-07 W=2e-06 AD=1.02e-12 AS=5.1e-13 PD=3.02e-06
+ PS=5.1e-07
mXI18.MM1 N_NET27_XI18.MM1_d N_A_XI18.MM1_g N_VDD_XI18.MM1_s N_VDD_XI20.MM0_b
+ P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI18.MM0 N_NET27_XI18.MM0_d N_CLKOUT_XI18.MM0_g N_VDD_XI18.MM0_s
+ N_VDD_XI20.MM0_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=5.1e-13 PD=5.1e-07
+ PS=2.02e-06
mXI20.MM1 N_NET25_XI20.MM1_d N_NET27_XI20.MM1_g N_VSS_XI20.MM1_s
+ N_VSS_XI20.MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI20.MM0 N_NET25_XI20.MM0_d N_NET27_XI20.MM0_g N_VDD_XI20.MM0_s
+ N_VDD_XI20.MM0_b P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06
+ PS=3.98e-06
mXI21.MM1 N_NET24_XI21.MM1_d N_NET25_XI21.MM1_g N_VSS_XI21.MM1_s
+ N_VSS_XI20.MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI21.MM0 N_NET24_XI21.MM0_d N_NET25_XI21.MM0_g N_VDD_XI21.MM0_s
+ N_VDD_XI20.MM0_b P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06
+ PS=3.98e-06
mXI22.MM1 N_NET23_XI22.MM1_d N_NET24_XI22.MM1_g N_VSS_XI22.MM1_s
+ N_VSS_XI20.MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI22.MM0 N_NET23_XI22.MM0_d N_NET24_XI22.MM0_g N_VDD_XI22.MM0_s
+ N_VDD_XI20.MM0_b P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06
+ PS=3.98e-06
mXI23.MM1 N_NET26_XI23.MM1_d N_NET23_XI23.MM1_g N_VSS_XI23.MM1_s
+ N_VSS_XI20.MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI23.MM0 N_NET26_XI23.MM0_d N_NET23_XI23.MM0_g N_VDD_XI23.MM0_s
+ N_VDD_XI20.MM0_b P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06
+ PS=3.98e-06
mXI24.MM1 N_NET023_XI24.MM1_d N_NET26_XI24.MM1_g N_VSS_XI24.MM1_s
+ N_VSS_XI20.MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI24.MM0 N_NET023_XI24.MM0_d N_NET26_XI24.MM0_g N_VDD_XI24.MM0_s
+ N_VDD_XI20.MM0_b P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06
+ PS=3.98e-06
mXI25.MM1 N_CLKOUT_XI25.MM1_d N_NET023_XI25.MM1_g N_VSS_XI25.MM1_s
+ N_VSS_XI20.MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI25.MM0 N_CLKOUT_XI25.MM0_d N_NET023_XI25.MM0_g N_VDD_XI25.MM0_s
+ N_VDD_XI20.MM0_b P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06
+ PS=3.98e-06
*
.include "/home/IC/lab6/CLKGEN/clkgen.pex.spi.CLKGEN.pxi"
*
.ends
*
*
