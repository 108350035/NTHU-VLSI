* File: /home/IC/final/READ/read_out.pex.spi
* Created: Thu Apr  3 17:16:18 2025
* Program "Calibre xRC"
* Version "v2019.3_15.11"
* 
.include "/home/IC/final/READ/read_out.pex.spi.pex"
.subckt read_out  EN RST CLK BL1 BL3 BL5 BL7 BL0 BL2 BL4 BL6 VSS VDD WL1 WL3 WL5
+ WL7 WL0 WL2 WL4 WL6
* 
* WL6	WL6
* WL4	WL4
* WL2	WL2
* WL0	WL0
* WL7	WL7
* WL5	WL5
* WL3	WL3
* WL1	WL1
* VDD	VDD
* VSS	VSS
* BL6	BL6
* BL4	BL4
* BL2	BL2
* BL0	BL0
* BL7	BL7
* BL5	BL5
* BL3	BL3
* BL1	BL1
* CLK	CLK
* RST	RST
* EN	EN
mXI1.XI52.MM14 N_BL1_XI1.XI52.MM14_d N_XI1.XI52.NET031_XI1.XI52.MM14_g
+ N_VSS_XI1.XI52.MM14_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI54.MM14 N_BL3_XI1.XI54.MM14_d N_XI1.XI54.NET031_XI1.XI54.MM14_g
+ N_VSS_XI1.XI54.MM14_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI56.MM14 N_BL5_XI1.XI56.MM14_d N_XI1.XI56.NET031_XI1.XI56.MM14_g
+ N_VSS_XI1.XI56.MM14_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI58.MM14 N_BL7_XI1.XI58.MM14_d N_XI1.XI58.NET031_XI1.XI58.MM14_g
+ N_VSS_XI1.XI58.MM14_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI52.MM14@4 N_BL1_XI1.XI52.MM14@4_d N_XI1.XI52.NET031_XI1.XI52.MM14@4_g
+ N_VSS_XI1.XI52.MM14@4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI54.MM14@4 N_BL3_XI1.XI54.MM14@4_d N_XI1.XI54.NET031_XI1.XI54.MM14@4_g
+ N_VSS_XI1.XI54.MM14@4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI56.MM14@4 N_BL5_XI1.XI56.MM14@4_d N_XI1.XI56.NET031_XI1.XI56.MM14@4_g
+ N_VSS_XI1.XI56.MM14@4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI58.MM14@4 N_BL7_XI1.XI58.MM14@4_d N_XI1.XI58.NET031_XI1.XI58.MM14@4_g
+ N_VSS_XI1.XI58.MM14@4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI52.MM14@3 N_BL1_XI1.XI52.MM14@3_d N_XI1.XI52.NET031_XI1.XI52.MM14@3_g
+ N_VSS_XI1.XI52.MM14@3_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI54.MM14@3 N_BL3_XI1.XI54.MM14@3_d N_XI1.XI54.NET031_XI1.XI54.MM14@3_g
+ N_VSS_XI1.XI54.MM14@3_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI56.MM14@3 N_BL5_XI1.XI56.MM14@3_d N_XI1.XI56.NET031_XI1.XI56.MM14@3_g
+ N_VSS_XI1.XI56.MM14@3_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI58.MM14@3 N_BL7_XI1.XI58.MM14@3_d N_XI1.XI58.NET031_XI1.XI58.MM14@3_g
+ N_VSS_XI1.XI58.MM14@3_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI52.MM14@2 N_BL1_XI1.XI52.MM14@2_d N_XI1.XI52.NET031_XI1.XI52.MM14@2_g
+ N_VSS_XI1.XI52.MM14@2_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI54.MM14@2 N_BL3_XI1.XI54.MM14@2_d N_XI1.XI54.NET031_XI1.XI54.MM14@2_g
+ N_VSS_XI1.XI54.MM14@2_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI56.MM14@2 N_BL5_XI1.XI56.MM14@2_d N_XI1.XI56.NET031_XI1.XI56.MM14@2_g
+ N_VSS_XI1.XI56.MM14@2_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI58.MM14@2 N_BL7_XI1.XI58.MM14@2_d N_XI1.XI58.NET031_XI1.XI58.MM14@2_g
+ N_VSS_XI1.XI58.MM14@2_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI52.MM13 N_XI1.XI52.NET031_XI1.XI52.MM13_d N_NET37_XI1.XI52.MM13_g
+ N_XI1.XI52.NET037_XI1.XI52.MM13_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07
+ AD=2.94e-13 AS=1.53e-13 PD=1.58e-06 PS=5.1e-07
mXI1.XI54.MM13 N_XI1.XI54.NET031_XI1.XI54.MM13_d N_NET37_XI1.XI54.MM13_g
+ N_XI1.XI54.NET037_XI1.XI54.MM13_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07
+ AD=2.94e-13 AS=1.53e-13 PD=1.58e-06 PS=5.1e-07
mXI1.XI56.MM13 N_XI1.XI56.NET031_XI1.XI56.MM13_d N_NET37_XI1.XI56.MM13_g
+ N_XI1.XI56.NET037_XI1.XI56.MM13_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07
+ AD=2.94e-13 AS=1.53e-13 PD=1.58e-06 PS=5.1e-07
mXI1.XI58.MM13 N_XI1.XI58.NET031_XI1.XI58.MM13_d N_NET37_XI1.XI58.MM13_g
+ N_XI1.XI58.NET037_XI1.XI58.MM13_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07
+ AD=2.94e-13 AS=1.53e-13 PD=1.58e-06 PS=5.1e-07
mXI1.XI52.MM12 N_XI1.XI52.NET037_XI1.XI52.MM12_d N_NET39_XI1.XI52.MM12_g
+ N_XI1.XI52.NET036_XI1.XI52.MM12_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07
+ AD=1.53e-13 AS=1.53e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI54.MM12 N_XI1.XI54.NET037_XI1.XI54.MM12_d N_NET41_XI1.XI54.MM12_g
+ N_XI1.XI54.NET036_XI1.XI54.MM12_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07
+ AD=1.53e-13 AS=1.53e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI56.MM12 N_XI1.XI56.NET037_XI1.XI56.MM12_d N_NET39_XI1.XI56.MM12_g
+ N_XI1.XI56.NET036_XI1.XI56.MM12_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07
+ AD=1.53e-13 AS=1.53e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI58.MM12 N_XI1.XI58.NET037_XI1.XI58.MM12_d N_NET41_XI1.XI58.MM12_g
+ N_XI1.XI58.NET036_XI1.XI58.MM12_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07
+ AD=1.53e-13 AS=1.53e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI52.MM11 N_XI1.XI52.NET036_XI1.XI52.MM11_d N_NET45_XI1.XI52.MM11_g
+ N_VSS_XI1.XI52.MM11_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07 AD=1.53e-13
+ AS=2.94e-13 PD=5.1e-07 PS=1.58e-06
mXI1.XI54.MM11 N_XI1.XI54.NET036_XI1.XI54.MM11_d N_NET45_XI1.XI54.MM11_g
+ N_VSS_XI1.XI54.MM11_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07 AD=1.53e-13
+ AS=2.94e-13 PD=5.1e-07 PS=1.58e-06
mXI1.XI56.MM11 N_XI1.XI56.NET036_XI1.XI56.MM11_d N_NET43_XI1.XI56.MM11_g
+ N_VSS_XI1.XI56.MM11_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07 AD=1.53e-13
+ AS=2.94e-13 PD=5.1e-07 PS=1.58e-06
mXI1.XI58.MM11 N_XI1.XI58.NET036_XI1.XI58.MM11_d N_NET43_XI1.XI58.MM11_g
+ N_VSS_XI1.XI58.MM11_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07 AD=1.53e-13
+ AS=2.94e-13 PD=5.1e-07 PS=1.58e-06
mXI1.XI43.MM11 N_XI1.XI43.NET036_XI1.XI43.MM11_d N_NET45_XI1.XI43.MM11_g
+ N_VSS_XI1.XI43.MM11_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07 AD=1.53e-13
+ AS=2.94e-13 PD=5.1e-07 PS=1.58e-06
mXI1.XI53.MM11 N_XI1.XI53.NET036_XI1.XI53.MM11_d N_NET45_XI1.XI53.MM11_g
+ N_VSS_XI1.XI53.MM11_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07 AD=1.53e-13
+ AS=2.94e-13 PD=5.1e-07 PS=1.58e-06
mXI1.XI55.MM11 N_XI1.XI55.NET036_XI1.XI55.MM11_d N_NET43_XI1.XI55.MM11_g
+ N_VSS_XI1.XI55.MM11_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07 AD=1.53e-13
+ AS=2.94e-13 PD=5.1e-07 PS=1.58e-06
mXI1.XI57.MM11 N_XI1.XI57.NET036_XI1.XI57.MM11_d N_NET43_XI1.XI57.MM11_g
+ N_VSS_XI1.XI57.MM11_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07 AD=1.53e-13
+ AS=2.94e-13 PD=5.1e-07 PS=1.58e-06
mXI1.XI43.MM12 N_XI1.XI43.NET037_XI1.XI43.MM12_d N_NET39_XI1.XI43.MM12_g
+ N_XI1.XI43.NET036_XI1.XI43.MM12_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07
+ AD=1.53e-13 AS=1.53e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI53.MM12 N_XI1.XI53.NET037_XI1.XI53.MM12_d N_NET41_XI1.XI53.MM12_g
+ N_XI1.XI53.NET036_XI1.XI53.MM12_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07
+ AD=1.53e-13 AS=1.53e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI55.MM12 N_XI1.XI55.NET037_XI1.XI55.MM12_d N_NET39_XI1.XI55.MM12_g
+ N_XI1.XI55.NET036_XI1.XI55.MM12_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07
+ AD=1.53e-13 AS=1.53e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI57.MM12 N_XI1.XI57.NET037_XI1.XI57.MM12_d N_NET41_XI1.XI57.MM12_g
+ N_XI1.XI57.NET036_XI1.XI57.MM12_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07
+ AD=1.53e-13 AS=1.53e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI43.MM13 N_XI1.XI43.NET031_XI1.XI43.MM13_d N_NET38_XI1.XI43.MM13_g
+ N_XI1.XI43.NET037_XI1.XI43.MM13_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07
+ AD=2.94e-13 AS=1.53e-13 PD=1.58e-06 PS=5.1e-07
mXI1.XI53.MM13 N_XI1.XI53.NET031_XI1.XI53.MM13_d N_NET38_XI1.XI53.MM13_g
+ N_XI1.XI53.NET037_XI1.XI53.MM13_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07
+ AD=2.94e-13 AS=1.53e-13 PD=1.58e-06 PS=5.1e-07
mXI1.XI55.MM13 N_XI1.XI55.NET031_XI1.XI55.MM13_d N_NET38_XI1.XI55.MM13_g
+ N_XI1.XI55.NET037_XI1.XI55.MM13_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07
+ AD=2.94e-13 AS=1.53e-13 PD=1.58e-06 PS=5.1e-07
mXI1.XI57.MM13 N_XI1.XI57.NET031_XI1.XI57.MM13_d N_NET38_XI1.XI57.MM13_g
+ N_XI1.XI57.NET037_XI1.XI57.MM13_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=6e-07
+ AD=2.94e-13 AS=1.53e-13 PD=1.58e-06 PS=5.1e-07
mXI1.XI43.MM14 N_BL0_XI1.XI43.MM14_d N_XI1.XI43.NET031_XI1.XI43.MM14_g
+ N_VSS_XI1.XI43.MM14_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI53.MM14 N_BL2_XI1.XI53.MM14_d N_XI1.XI53.NET031_XI1.XI53.MM14_g
+ N_VSS_XI1.XI53.MM14_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI55.MM14 N_BL4_XI1.XI55.MM14_d N_XI1.XI55.NET031_XI1.XI55.MM14_g
+ N_VSS_XI1.XI55.MM14_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI57.MM14 N_BL6_XI1.XI57.MM14_d N_XI1.XI57.NET031_XI1.XI57.MM14_g
+ N_VSS_XI1.XI57.MM14_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI43.MM14@4 N_BL0_XI1.XI43.MM14@4_d N_XI1.XI43.NET031_XI1.XI43.MM14@4_g
+ N_VSS_XI1.XI43.MM14@4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI53.MM14@4 N_BL2_XI1.XI53.MM14@4_d N_XI1.XI53.NET031_XI1.XI53.MM14@4_g
+ N_VSS_XI1.XI53.MM14@4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI55.MM14@4 N_BL4_XI1.XI55.MM14@4_d N_XI1.XI55.NET031_XI1.XI55.MM14@4_g
+ N_VSS_XI1.XI55.MM14@4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI57.MM14@4 N_BL6_XI1.XI57.MM14@4_d N_XI1.XI57.NET031_XI1.XI57.MM14@4_g
+ N_VSS_XI1.XI57.MM14@4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI43.MM14@3 N_BL0_XI1.XI43.MM14@3_d N_XI1.XI43.NET031_XI1.XI43.MM14@3_g
+ N_VSS_XI1.XI43.MM14@3_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI53.MM14@3 N_BL2_XI1.XI53.MM14@3_d N_XI1.XI53.NET031_XI1.XI53.MM14@3_g
+ N_VSS_XI1.XI53.MM14@3_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI55.MM14@3 N_BL4_XI1.XI55.MM14@3_d N_XI1.XI55.NET031_XI1.XI55.MM14@3_g
+ N_VSS_XI1.XI55.MM14@3_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI57.MM14@3 N_BL6_XI1.XI57.MM14@3_d N_XI1.XI57.NET031_XI1.XI57.MM14@3_g
+ N_VSS_XI1.XI57.MM14@3_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI43.MM14@2 N_BL0_XI1.XI43.MM14@2_d N_XI1.XI43.NET031_XI1.XI43.MM14@2_g
+ N_VSS_XI1.XI43.MM14@2_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI53.MM14@2 N_BL2_XI1.XI53.MM14@2_d N_XI1.XI53.NET031_XI1.XI53.MM14@2_g
+ N_VSS_XI1.XI53.MM14@2_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI55.MM14@2 N_BL4_XI1.XI55.MM14@2_d N_XI1.XI55.NET031_XI1.XI55.MM14@2_g
+ N_VSS_XI1.XI55.MM14@2_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI57.MM14@2 N_BL6_XI1.XI57.MM14@2_d N_XI1.XI57.NET031_XI1.XI57.MM14@2_g
+ N_VSS_XI1.XI57.MM14@2_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI52.MM14 N_WL1_XI2.XI52.MM14_d N_XI2.XI52.NET031_XI2.XI52.MM14_g
+ N_VSS_XI2.XI52.MM14_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI54.MM14 N_WL3_XI2.XI54.MM14_d N_XI2.XI54.NET031_XI2.XI54.MM14_g
+ N_VSS_XI2.XI54.MM14_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI56.MM14 N_WL5_XI2.XI56.MM14_d N_XI2.XI56.NET031_XI2.XI56.MM14_g
+ N_VSS_XI2.XI56.MM14_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI58.MM14 N_WL7_XI2.XI58.MM14_d N_XI2.XI58.NET031_XI2.XI58.MM14_g
+ N_VSS_XI2.XI58.MM14_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI52.MM14@4 N_WL1_XI2.XI52.MM14@4_d N_XI2.XI52.NET031_XI2.XI52.MM14@4_g
+ N_VSS_XI2.XI52.MM14@4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI54.MM14@4 N_WL3_XI2.XI54.MM14@4_d N_XI2.XI54.NET031_XI2.XI54.MM14@4_g
+ N_VSS_XI2.XI54.MM14@4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI56.MM14@4 N_WL5_XI2.XI56.MM14@4_d N_XI2.XI56.NET031_XI2.XI56.MM14@4_g
+ N_VSS_XI2.XI56.MM14@4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI58.MM14@4 N_WL7_XI2.XI58.MM14@4_d N_XI2.XI58.NET031_XI2.XI58.MM14@4_g
+ N_VSS_XI2.XI58.MM14@4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI52.MM14@3 N_WL1_XI2.XI52.MM14@3_d N_XI2.XI52.NET031_XI2.XI52.MM14@3_g
+ N_VSS_XI2.XI52.MM14@3_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI54.MM14@3 N_WL3_XI2.XI54.MM14@3_d N_XI2.XI54.NET031_XI2.XI54.MM14@3_g
+ N_VSS_XI2.XI54.MM14@3_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI56.MM14@3 N_WL5_XI2.XI56.MM14@3_d N_XI2.XI56.NET031_XI2.XI56.MM14@3_g
+ N_VSS_XI2.XI56.MM14@3_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI58.MM14@3 N_WL7_XI2.XI58.MM14@3_d N_XI2.XI58.NET031_XI2.XI58.MM14@3_g
+ N_VSS_XI2.XI58.MM14@3_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI52.MM14@2 N_WL1_XI2.XI52.MM14@2_d N_XI2.XI52.NET031_XI2.XI52.MM14@2_g
+ N_VSS_XI2.XI52.MM14@2_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI54.MM14@2 N_WL3_XI2.XI54.MM14@2_d N_XI2.XI54.NET031_XI2.XI54.MM14@2_g
+ N_VSS_XI2.XI54.MM14@2_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI56.MM14@2 N_WL5_XI2.XI56.MM14@2_d N_XI2.XI56.NET031_XI2.XI56.MM14@2_g
+ N_VSS_XI2.XI56.MM14@2_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI58.MM14@2 N_WL7_XI2.XI58.MM14@2_d N_XI2.XI58.NET031_XI2.XI58.MM14@2_g
+ N_VSS_XI2.XI58.MM14@2_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI52.MM13 N_XI2.XI52.NET031_XI2.XI52.MM13_d N_NET47_XI2.XI52.MM13_g
+ N_XI2.XI52.NET036_XI2.XI52.MM13_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI2.XI54.MM13 N_XI2.XI54.NET031_XI2.XI54.MM13_d N_NET47_XI2.XI54.MM13_g
+ N_XI2.XI54.NET036_XI2.XI54.MM13_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI2.XI56.MM13 N_XI2.XI56.NET031_XI2.XI56.MM13_d N_NET47_XI2.XI56.MM13_g
+ N_XI2.XI56.NET036_XI2.XI56.MM13_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI2.XI58.MM13 N_XI2.XI58.NET031_XI2.XI58.MM13_d N_NET47_XI2.XI58.MM13_g
+ N_XI2.XI58.NET036_XI2.XI58.MM13_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI2.XI52.MM12 N_XI2.XI52.NET036_XI2.XI52.MM12_d N_NET44_XI2.XI52.MM12_g
+ N_XI2.XI52.NET037_XI2.XI52.MM12_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI54.MM12 N_XI2.XI54.NET036_XI2.XI54.MM12_d N_NET46_XI2.XI54.MM12_g
+ N_XI2.XI54.NET037_XI2.XI54.MM12_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI56.MM12 N_XI2.XI56.NET036_XI2.XI56.MM12_d N_NET44_XI2.XI56.MM12_g
+ N_XI2.XI56.NET037_XI2.XI56.MM12_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI58.MM12 N_XI2.XI58.NET036_XI2.XI58.MM12_d N_NET46_XI2.XI58.MM12_g
+ N_XI2.XI58.NET037_XI2.XI58.MM12_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI52.MM11 N_XI2.XI52.NET037_XI2.XI52.MM11_d N_NET40_XI2.XI52.MM11_g
+ N_VSS_XI2.XI52.MM11_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI2.XI54.MM11 N_XI2.XI54.NET037_XI2.XI54.MM11_d N_NET40_XI2.XI54.MM11_g
+ N_VSS_XI2.XI54.MM11_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI2.XI56.MM11 N_XI2.XI56.NET037_XI2.XI56.MM11_d N_NET42_XI2.XI56.MM11_g
+ N_VSS_XI2.XI56.MM11_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI2.XI58.MM11 N_XI2.XI58.NET037_XI2.XI58.MM11_d N_NET42_XI2.XI58.MM11_g
+ N_VSS_XI2.XI58.MM11_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI2.XI43.MM11 N_XI2.XI43.NET037_XI2.XI43.MM11_d N_NET40_XI2.XI43.MM11_g
+ N_VSS_XI2.XI43.MM11_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI2.XI53.MM11 N_XI2.XI53.NET037_XI2.XI53.MM11_d N_NET40_XI2.XI53.MM11_g
+ N_VSS_XI2.XI53.MM11_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI2.XI55.MM11 N_XI2.XI55.NET037_XI2.XI55.MM11_d N_NET42_XI2.XI55.MM11_g
+ N_VSS_XI2.XI55.MM11_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI2.XI57.MM11 N_XI2.XI57.NET037_XI2.XI57.MM11_d N_NET42_XI2.XI57.MM11_g
+ N_VSS_XI2.XI57.MM11_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI2.XI43.MM12 N_XI2.XI43.NET036_XI2.XI43.MM12_d N_NET44_XI2.XI43.MM12_g
+ N_XI2.XI43.NET037_XI2.XI43.MM12_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI53.MM12 N_XI2.XI53.NET036_XI2.XI53.MM12_d N_NET46_XI2.XI53.MM12_g
+ N_XI2.XI53.NET037_XI2.XI53.MM12_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI55.MM12 N_XI2.XI55.NET036_XI2.XI55.MM12_d N_NET44_XI2.XI55.MM12_g
+ N_XI2.XI55.NET037_XI2.XI55.MM12_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI57.MM12 N_XI2.XI57.NET036_XI2.XI57.MM12_d N_NET46_XI2.XI57.MM12_g
+ N_XI2.XI57.NET037_XI2.XI57.MM12_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI43.MM13 N_XI2.XI43.NET031_XI2.XI43.MM13_d N_NET48_XI2.XI43.MM13_g
+ N_XI2.XI43.NET036_XI2.XI43.MM13_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI2.XI53.MM13 N_XI2.XI53.NET031_XI2.XI53.MM13_d N_NET48_XI2.XI53.MM13_g
+ N_XI2.XI53.NET036_XI2.XI53.MM13_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI2.XI55.MM13 N_XI2.XI55.NET031_XI2.XI55.MM13_d N_NET48_XI2.XI55.MM13_g
+ N_XI2.XI55.NET036_XI2.XI55.MM13_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI2.XI57.MM13 N_XI2.XI57.NET031_XI2.XI57.MM13_d N_NET48_XI2.XI57.MM13_g
+ N_XI2.XI57.NET036_XI2.XI57.MM13_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI2.XI43.MM14 N_WL0_XI2.XI43.MM14_d N_XI2.XI43.NET031_XI2.XI43.MM14_g
+ N_VSS_XI2.XI43.MM14_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI53.MM14 N_WL2_XI2.XI53.MM14_d N_XI2.XI53.NET031_XI2.XI53.MM14_g
+ N_VSS_XI2.XI53.MM14_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI55.MM14 N_WL4_XI2.XI55.MM14_d N_XI2.XI55.NET031_XI2.XI55.MM14_g
+ N_VSS_XI2.XI55.MM14_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI57.MM14 N_WL6_XI2.XI57.MM14_d N_XI2.XI57.NET031_XI2.XI57.MM14_g
+ N_VSS_XI2.XI57.MM14_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI43.MM14@4 N_WL0_XI2.XI43.MM14@4_d N_XI2.XI43.NET031_XI2.XI43.MM14@4_g
+ N_VSS_XI2.XI43.MM14@4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI53.MM14@4 N_WL2_XI2.XI53.MM14@4_d N_XI2.XI53.NET031_XI2.XI53.MM14@4_g
+ N_VSS_XI2.XI53.MM14@4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI55.MM14@4 N_WL4_XI2.XI55.MM14@4_d N_XI2.XI55.NET031_XI2.XI55.MM14@4_g
+ N_VSS_XI2.XI55.MM14@4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI57.MM14@4 N_WL6_XI2.XI57.MM14@4_d N_XI2.XI57.NET031_XI2.XI57.MM14@4_g
+ N_VSS_XI2.XI57.MM14@4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI43.MM14@3 N_WL0_XI2.XI43.MM14@3_d N_XI2.XI43.NET031_XI2.XI43.MM14@3_g
+ N_VSS_XI2.XI43.MM14@3_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI53.MM14@3 N_WL2_XI2.XI53.MM14@3_d N_XI2.XI53.NET031_XI2.XI53.MM14@3_g
+ N_VSS_XI2.XI53.MM14@3_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI55.MM14@3 N_WL4_XI2.XI55.MM14@3_d N_XI2.XI55.NET031_XI2.XI55.MM14@3_g
+ N_VSS_XI2.XI55.MM14@3_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI57.MM14@3 N_WL6_XI2.XI57.MM14@3_d N_XI2.XI57.NET031_XI2.XI57.MM14@3_g
+ N_VSS_XI2.XI57.MM14@3_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI43.MM14@2 N_WL0_XI2.XI43.MM14@2_d N_XI2.XI43.NET031_XI2.XI43.MM14@2_g
+ N_VSS_XI2.XI43.MM14@2_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI53.MM14@2 N_WL2_XI2.XI53.MM14@2_d N_XI2.XI53.NET031_XI2.XI53.MM14@2_g
+ N_VSS_XI2.XI53.MM14@2_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI55.MM14@2 N_WL4_XI2.XI55.MM14@2_d N_XI2.XI55.NET031_XI2.XI55.MM14@2_g
+ N_VSS_XI2.XI55.MM14@2_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI57.MM14@2 N_WL6_XI2.XI57.MM14@2_d N_XI2.XI57.NET031_XI2.XI57.MM14@2_g
+ N_VSS_XI2.XI57.MM14@2_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI52.MM18 N_BL1_XI1.XI52.MM18_d N_XI1.XI52.NET031_XI1.XI52.MM18_g
+ N_VDD_XI1.XI52.MM18_s N_VDD_XI1.XI52.MM18_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI54.MM18 N_BL3_XI1.XI54.MM18_d N_XI1.XI54.NET031_XI1.XI54.MM18_g
+ N_VDD_XI1.XI54.MM18_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI56.MM18 N_BL5_XI1.XI56.MM18_d N_XI1.XI56.NET031_XI1.XI56.MM18_g
+ N_VDD_XI1.XI56.MM18_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI58.MM18 N_BL7_XI1.XI58.MM18_d N_XI1.XI58.NET031_XI1.XI58.MM18_g
+ N_VDD_XI1.XI58.MM18_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI52.MM18@4 N_BL1_XI1.XI52.MM18@4_d N_XI1.XI52.NET031_XI1.XI52.MM18@4_g
+ N_VDD_XI1.XI52.MM18@4_s N_VDD_XI1.XI52.MM18_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI54.MM18@4 N_BL3_XI1.XI54.MM18@4_d N_XI1.XI54.NET031_XI1.XI54.MM18@4_g
+ N_VDD_XI1.XI54.MM18@4_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI56.MM18@4 N_BL5_XI1.XI56.MM18@4_d N_XI1.XI56.NET031_XI1.XI56.MM18@4_g
+ N_VDD_XI1.XI56.MM18@4_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI58.MM18@4 N_BL7_XI1.XI58.MM18@4_d N_XI1.XI58.NET031_XI1.XI58.MM18@4_g
+ N_VDD_XI1.XI58.MM18@4_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI52.MM18@3 N_BL1_XI1.XI52.MM18@3_d N_XI1.XI52.NET031_XI1.XI52.MM18@3_g
+ N_VDD_XI1.XI52.MM18@3_s N_VDD_XI1.XI52.MM18_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI54.MM18@3 N_BL3_XI1.XI54.MM18@3_d N_XI1.XI54.NET031_XI1.XI54.MM18@3_g
+ N_VDD_XI1.XI54.MM18@3_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI56.MM18@3 N_BL5_XI1.XI56.MM18@3_d N_XI1.XI56.NET031_XI1.XI56.MM18@3_g
+ N_VDD_XI1.XI56.MM18@3_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI58.MM18@3 N_BL7_XI1.XI58.MM18@3_d N_XI1.XI58.NET031_XI1.XI58.MM18@3_g
+ N_VDD_XI1.XI58.MM18@3_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI52.MM18@2 N_BL1_XI1.XI52.MM18@2_d N_XI1.XI52.NET031_XI1.XI52.MM18@2_g
+ N_VDD_XI1.XI52.MM18@2_s N_VDD_XI1.XI52.MM18_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI54.MM18@2 N_BL3_XI1.XI54.MM18@2_d N_XI1.XI54.NET031_XI1.XI54.MM18@2_g
+ N_VDD_XI1.XI54.MM18@2_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI56.MM18@2 N_BL5_XI1.XI56.MM18@2_d N_XI1.XI56.NET031_XI1.XI56.MM18@2_g
+ N_VDD_XI1.XI56.MM18@2_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI58.MM18@2 N_BL7_XI1.XI58.MM18@2_d N_XI1.XI58.NET031_XI1.XI58.MM18@2_g
+ N_VDD_XI1.XI58.MM18@2_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI52.MM17 N_XI1.XI52.NET031_XI1.XI52.MM17_d N_EN_XI1.XI52.MM17_g
+ N_VDD_XI1.XI52.MM17_s N_VDD_XI1.XI52.MM18_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI1.XI54.MM17 N_XI1.XI54.NET031_XI1.XI54.MM17_d N_EN_XI1.XI54.MM17_g
+ N_VDD_XI1.XI54.MM17_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI1.XI56.MM17 N_XI1.XI56.NET031_XI1.XI56.MM17_d N_EN_XI1.XI56.MM17_g
+ N_VDD_XI1.XI56.MM17_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI1.XI58.MM17 N_XI1.XI58.NET031_XI1.XI58.MM17_d N_EN_XI1.XI58.MM17_g
+ N_VDD_XI1.XI58.MM17_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI1.XI52.MM15 N_XI1.XI52.NET031_XI1.XI52.MM15_d N_NET37_XI1.XI52.MM15_g
+ N_VDD_XI1.XI52.MM15_s N_VDD_XI1.XI52.MM18_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI54.MM15 N_XI1.XI54.NET031_XI1.XI54.MM15_d N_NET37_XI1.XI54.MM15_g
+ N_VDD_XI1.XI54.MM15_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI56.MM15 N_XI1.XI56.NET031_XI1.XI56.MM15_d N_NET37_XI1.XI56.MM15_g
+ N_VDD_XI1.XI56.MM15_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI58.MM15 N_XI1.XI58.NET031_XI1.XI58.MM15_d N_NET37_XI1.XI58.MM15_g
+ N_VDD_XI1.XI58.MM15_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI52.MM16 N_XI1.XI52.NET031_XI1.XI52.MM16_d N_NET39_XI1.XI52.MM16_g
+ N_VDD_XI1.XI52.MM16_s N_VDD_XI1.XI52.MM18_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI54.MM16 N_XI1.XI54.NET031_XI1.XI54.MM16_d N_NET41_XI1.XI54.MM16_g
+ N_VDD_XI1.XI54.MM16_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI56.MM16 N_XI1.XI56.NET031_XI1.XI56.MM16_d N_NET39_XI1.XI56.MM16_g
+ N_VDD_XI1.XI56.MM16_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI58.MM16 N_XI1.XI58.NET031_XI1.XI58.MM16_d N_NET41_XI1.XI58.MM16_g
+ N_VDD_XI1.XI58.MM16_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI52.MM19 N_XI1.XI52.NET031_XI1.XI52.MM19_d N_NET45_XI1.XI52.MM19_g
+ N_VDD_XI1.XI52.MM19_s N_VDD_XI1.XI52.MM18_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI1.XI54.MM19 N_XI1.XI54.NET031_XI1.XI54.MM19_d N_NET45_XI1.XI54.MM19_g
+ N_VDD_XI1.XI54.MM19_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI1.XI56.MM19 N_XI1.XI56.NET031_XI1.XI56.MM19_d N_NET43_XI1.XI56.MM19_g
+ N_VDD_XI1.XI56.MM19_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI1.XI58.MM19 N_XI1.XI58.NET031_XI1.XI58.MM19_d N_NET43_XI1.XI58.MM19_g
+ N_VDD_XI1.XI58.MM19_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI1.XI43.MM19 N_XI1.XI43.NET031_XI1.XI43.MM19_d N_NET45_XI1.XI43.MM19_g
+ N_VDD_XI1.XI43.MM19_s N_VDD_XI1.XI52.MM18_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI1.XI53.MM19 N_XI1.XI53.NET031_XI1.XI53.MM19_d N_NET45_XI1.XI53.MM19_g
+ N_VDD_XI1.XI53.MM19_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI1.XI55.MM19 N_XI1.XI55.NET031_XI1.XI55.MM19_d N_NET43_XI1.XI55.MM19_g
+ N_VDD_XI1.XI55.MM19_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI1.XI57.MM19 N_XI1.XI57.NET031_XI1.XI57.MM19_d N_NET43_XI1.XI57.MM19_g
+ N_VDD_XI1.XI57.MM19_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI1.XI43.MM16 N_XI1.XI43.NET031_XI1.XI43.MM16_d N_NET39_XI1.XI43.MM16_g
+ N_VDD_XI1.XI43.MM16_s N_VDD_XI1.XI52.MM18_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI53.MM16 N_XI1.XI53.NET031_XI1.XI53.MM16_d N_NET41_XI1.XI53.MM16_g
+ N_VDD_XI1.XI53.MM16_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI55.MM16 N_XI1.XI55.NET031_XI1.XI55.MM16_d N_NET39_XI1.XI55.MM16_g
+ N_VDD_XI1.XI55.MM16_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI57.MM16 N_XI1.XI57.NET031_XI1.XI57.MM16_d N_NET41_XI1.XI57.MM16_g
+ N_VDD_XI1.XI57.MM16_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI43.MM15 N_XI1.XI43.NET031_XI1.XI43.MM15_d N_NET38_XI1.XI43.MM15_g
+ N_VDD_XI1.XI43.MM15_s N_VDD_XI1.XI52.MM18_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI53.MM15 N_XI1.XI53.NET031_XI1.XI53.MM15_d N_NET38_XI1.XI53.MM15_g
+ N_VDD_XI1.XI53.MM15_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI55.MM15 N_XI1.XI55.NET031_XI1.XI55.MM15_d N_NET38_XI1.XI55.MM15_g
+ N_VDD_XI1.XI55.MM15_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI57.MM15 N_XI1.XI57.NET031_XI1.XI57.MM15_d N_NET38_XI1.XI57.MM15_g
+ N_VDD_XI1.XI57.MM15_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI43.MM17 N_XI1.XI43.NET031_XI1.XI43.MM17_d N_EN_XI1.XI43.MM17_g
+ N_VDD_XI1.XI43.MM17_s N_VDD_XI1.XI52.MM18_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI1.XI53.MM17 N_XI1.XI53.NET031_XI1.XI53.MM17_d N_EN_XI1.XI53.MM17_g
+ N_VDD_XI1.XI53.MM17_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI1.XI55.MM17 N_XI1.XI55.NET031_XI1.XI55.MM17_d N_EN_XI1.XI55.MM17_g
+ N_VDD_XI1.XI55.MM17_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI1.XI57.MM17 N_XI1.XI57.NET031_XI1.XI57.MM17_d N_EN_XI1.XI57.MM17_g
+ N_VDD_XI1.XI57.MM17_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI1.XI43.MM18 N_BL0_XI1.XI43.MM18_d N_XI1.XI43.NET031_XI1.XI43.MM18_g
+ N_VDD_XI1.XI43.MM18_s N_VDD_XI1.XI52.MM18_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI53.MM18 N_BL2_XI1.XI53.MM18_d N_XI1.XI53.NET031_XI1.XI53.MM18_g
+ N_VDD_XI1.XI53.MM18_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI55.MM18 N_BL4_XI1.XI55.MM18_d N_XI1.XI55.NET031_XI1.XI55.MM18_g
+ N_VDD_XI1.XI55.MM18_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI57.MM18 N_BL6_XI1.XI57.MM18_d N_XI1.XI57.NET031_XI1.XI57.MM18_g
+ N_VDD_XI1.XI57.MM18_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI43.MM18@4 N_BL0_XI1.XI43.MM18@4_d N_XI1.XI43.NET031_XI1.XI43.MM18@4_g
+ N_VDD_XI1.XI43.MM18@4_s N_VDD_XI1.XI52.MM18_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI53.MM18@4 N_BL2_XI1.XI53.MM18@4_d N_XI1.XI53.NET031_XI1.XI53.MM18@4_g
+ N_VDD_XI1.XI53.MM18@4_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI55.MM18@4 N_BL4_XI1.XI55.MM18@4_d N_XI1.XI55.NET031_XI1.XI55.MM18@4_g
+ N_VDD_XI1.XI55.MM18@4_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI57.MM18@4 N_BL6_XI1.XI57.MM18@4_d N_XI1.XI57.NET031_XI1.XI57.MM18@4_g
+ N_VDD_XI1.XI57.MM18@4_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI43.MM18@3 N_BL0_XI1.XI43.MM18@3_d N_XI1.XI43.NET031_XI1.XI43.MM18@3_g
+ N_VDD_XI1.XI43.MM18@3_s N_VDD_XI1.XI52.MM18_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI53.MM18@3 N_BL2_XI1.XI53.MM18@3_d N_XI1.XI53.NET031_XI1.XI53.MM18@3_g
+ N_VDD_XI1.XI53.MM18@3_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI55.MM18@3 N_BL4_XI1.XI55.MM18@3_d N_XI1.XI55.NET031_XI1.XI55.MM18@3_g
+ N_VDD_XI1.XI55.MM18@3_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI57.MM18@3 N_BL6_XI1.XI57.MM18@3_d N_XI1.XI57.NET031_XI1.XI57.MM18@3_g
+ N_VDD_XI1.XI57.MM18@3_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI43.MM18@2 N_BL0_XI1.XI43.MM18@2_d N_XI1.XI43.NET031_XI1.XI43.MM18@2_g
+ N_VDD_XI1.XI43.MM18@2_s N_VDD_XI1.XI52.MM18_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI53.MM18@2 N_BL2_XI1.XI53.MM18@2_d N_XI1.XI53.NET031_XI1.XI53.MM18@2_g
+ N_VDD_XI1.XI53.MM18@2_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI55.MM18@2 N_BL4_XI1.XI55.MM18@2_d N_XI1.XI55.NET031_XI1.XI55.MM18@2_g
+ N_VDD_XI1.XI55.MM18@2_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI57.MM18@2 N_BL6_XI1.XI57.MM18@2_d N_XI1.XI57.NET031_XI1.XI57.MM18@2_g
+ N_VDD_XI1.XI57.MM18@2_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI52.MM18 N_WL1_XI2.XI52.MM18_d N_XI2.XI52.NET031_XI2.XI52.MM18_g
+ N_VDD_XI2.XI52.MM18_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI54.MM18 N_WL3_XI2.XI54.MM18_d N_XI2.XI54.NET031_XI2.XI54.MM18_g
+ N_VDD_XI2.XI54.MM18_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI56.MM18 N_WL5_XI2.XI56.MM18_d N_XI2.XI56.NET031_XI2.XI56.MM18_g
+ N_VDD_XI2.XI56.MM18_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI58.MM18 N_WL7_XI2.XI58.MM18_d N_XI2.XI58.NET031_XI2.XI58.MM18_g
+ N_VDD_XI2.XI58.MM18_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI52.MM18@4 N_WL1_XI2.XI52.MM18@4_d N_XI2.XI52.NET031_XI2.XI52.MM18@4_g
+ N_VDD_XI2.XI52.MM18@4_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI54.MM18@4 N_WL3_XI2.XI54.MM18@4_d N_XI2.XI54.NET031_XI2.XI54.MM18@4_g
+ N_VDD_XI2.XI54.MM18@4_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI56.MM18@4 N_WL5_XI2.XI56.MM18@4_d N_XI2.XI56.NET031_XI2.XI56.MM18@4_g
+ N_VDD_XI2.XI56.MM18@4_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI58.MM18@4 N_WL7_XI2.XI58.MM18@4_d N_XI2.XI58.NET031_XI2.XI58.MM18@4_g
+ N_VDD_XI2.XI58.MM18@4_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI52.MM18@3 N_WL1_XI2.XI52.MM18@3_d N_XI2.XI52.NET031_XI2.XI52.MM18@3_g
+ N_VDD_XI2.XI52.MM18@3_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI54.MM18@3 N_WL3_XI2.XI54.MM18@3_d N_XI2.XI54.NET031_XI2.XI54.MM18@3_g
+ N_VDD_XI2.XI54.MM18@3_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI56.MM18@3 N_WL5_XI2.XI56.MM18@3_d N_XI2.XI56.NET031_XI2.XI56.MM18@3_g
+ N_VDD_XI2.XI56.MM18@3_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI58.MM18@3 N_WL7_XI2.XI58.MM18@3_d N_XI2.XI58.NET031_XI2.XI58.MM18@3_g
+ N_VDD_XI2.XI58.MM18@3_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI52.MM18@2 N_WL1_XI2.XI52.MM18@2_d N_XI2.XI52.NET031_XI2.XI52.MM18@2_g
+ N_VDD_XI2.XI52.MM18@2_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI54.MM18@2 N_WL3_XI2.XI54.MM18@2_d N_XI2.XI54.NET031_XI2.XI54.MM18@2_g
+ N_VDD_XI2.XI54.MM18@2_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI56.MM18@2 N_WL5_XI2.XI56.MM18@2_d N_XI2.XI56.NET031_XI2.XI56.MM18@2_g
+ N_VDD_XI2.XI56.MM18@2_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI58.MM18@2 N_WL7_XI2.XI58.MM18@2_d N_XI2.XI58.NET031_XI2.XI58.MM18@2_g
+ N_VDD_XI2.XI58.MM18@2_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI52.MM17 N_XI2.XI52.NET031_XI2.XI52.MM17_d N_EN_XI2.XI52.MM17_g
+ N_VDD_XI2.XI52.MM17_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI2.XI54.MM17 N_XI2.XI54.NET031_XI2.XI54.MM17_d N_EN_XI2.XI54.MM17_g
+ N_VDD_XI2.XI54.MM17_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI2.XI56.MM17 N_XI2.XI56.NET031_XI2.XI56.MM17_d N_EN_XI2.XI56.MM17_g
+ N_VDD_XI2.XI56.MM17_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI2.XI58.MM17 N_XI2.XI58.NET031_XI2.XI58.MM17_d N_EN_XI2.XI58.MM17_g
+ N_VDD_XI2.XI58.MM17_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI2.XI52.MM15 N_XI2.XI52.NET031_XI2.XI52.MM15_d N_NET47_XI2.XI52.MM15_g
+ N_VDD_XI2.XI52.MM15_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI54.MM15 N_XI2.XI54.NET031_XI2.XI54.MM15_d N_NET47_XI2.XI54.MM15_g
+ N_VDD_XI2.XI54.MM15_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI56.MM15 N_XI2.XI56.NET031_XI2.XI56.MM15_d N_NET47_XI2.XI56.MM15_g
+ N_VDD_XI2.XI56.MM15_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI58.MM15 N_XI2.XI58.NET031_XI2.XI58.MM15_d N_NET47_XI2.XI58.MM15_g
+ N_VDD_XI2.XI58.MM15_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI52.MM16 N_XI2.XI52.NET031_XI2.XI52.MM16_d N_NET44_XI2.XI52.MM16_g
+ N_VDD_XI2.XI52.MM16_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI54.MM16 N_XI2.XI54.NET031_XI2.XI54.MM16_d N_NET46_XI2.XI54.MM16_g
+ N_VDD_XI2.XI54.MM16_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI56.MM16 N_XI2.XI56.NET031_XI2.XI56.MM16_d N_NET44_XI2.XI56.MM16_g
+ N_VDD_XI2.XI56.MM16_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI58.MM16 N_XI2.XI58.NET031_XI2.XI58.MM16_d N_NET46_XI2.XI58.MM16_g
+ N_VDD_XI2.XI58.MM16_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI52.MM19 N_XI2.XI52.NET031_XI2.XI52.MM19_d N_NET40_XI2.XI52.MM19_g
+ N_VDD_XI2.XI52.MM19_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI2.XI54.MM19 N_XI2.XI54.NET031_XI2.XI54.MM19_d N_NET40_XI2.XI54.MM19_g
+ N_VDD_XI2.XI54.MM19_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI2.XI56.MM19 N_XI2.XI56.NET031_XI2.XI56.MM19_d N_NET42_XI2.XI56.MM19_g
+ N_VDD_XI2.XI56.MM19_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI2.XI58.MM19 N_XI2.XI58.NET031_XI2.XI58.MM19_d N_NET42_XI2.XI58.MM19_g
+ N_VDD_XI2.XI58.MM19_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI2.XI43.MM19 N_XI2.XI43.NET031_XI2.XI43.MM19_d N_NET40_XI2.XI43.MM19_g
+ N_VDD_XI2.XI43.MM19_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI2.XI53.MM19 N_XI2.XI53.NET031_XI2.XI53.MM19_d N_NET40_XI2.XI53.MM19_g
+ N_VDD_XI2.XI53.MM19_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI2.XI55.MM19 N_XI2.XI55.NET031_XI2.XI55.MM19_d N_NET42_XI2.XI55.MM19_g
+ N_VDD_XI2.XI55.MM19_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI2.XI57.MM19 N_XI2.XI57.NET031_XI2.XI57.MM19_d N_NET42_XI2.XI57.MM19_g
+ N_VDD_XI2.XI57.MM19_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI2.XI43.MM16 N_XI2.XI43.NET031_XI2.XI43.MM16_d N_NET44_XI2.XI43.MM16_g
+ N_VDD_XI2.XI43.MM16_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI53.MM16 N_XI2.XI53.NET031_XI2.XI53.MM16_d N_NET46_XI2.XI53.MM16_g
+ N_VDD_XI2.XI53.MM16_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI55.MM16 N_XI2.XI55.NET031_XI2.XI55.MM16_d N_NET44_XI2.XI55.MM16_g
+ N_VDD_XI2.XI55.MM16_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI57.MM16 N_XI2.XI57.NET031_XI2.XI57.MM16_d N_NET46_XI2.XI57.MM16_g
+ N_VDD_XI2.XI57.MM16_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI43.MM15 N_XI2.XI43.NET031_XI2.XI43.MM15_d N_NET48_XI2.XI43.MM15_g
+ N_VDD_XI2.XI43.MM15_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI53.MM15 N_XI2.XI53.NET031_XI2.XI53.MM15_d N_NET48_XI2.XI53.MM15_g
+ N_VDD_XI2.XI53.MM15_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI55.MM15 N_XI2.XI55.NET031_XI2.XI55.MM15_d N_NET48_XI2.XI55.MM15_g
+ N_VDD_XI2.XI55.MM15_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI57.MM15 N_XI2.XI57.NET031_XI2.XI57.MM15_d N_NET48_XI2.XI57.MM15_g
+ N_VDD_XI2.XI57.MM15_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI43.MM17 N_XI2.XI43.NET031_XI2.XI43.MM17_d N_EN_XI2.XI43.MM17_g
+ N_VDD_XI2.XI43.MM17_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI2.XI53.MM17 N_XI2.XI53.NET031_XI2.XI53.MM17_d N_EN_XI2.XI53.MM17_g
+ N_VDD_XI2.XI53.MM17_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI2.XI55.MM17 N_XI2.XI55.NET031_XI2.XI55.MM17_d N_EN_XI2.XI55.MM17_g
+ N_VDD_XI2.XI55.MM17_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI2.XI57.MM17 N_XI2.XI57.NET031_XI2.XI57.MM17_d N_EN_XI2.XI57.MM17_g
+ N_VDD_XI2.XI57.MM17_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=3.06e-13 PD=2.18e-06 PS=5.1e-07
mXI2.XI43.MM18 N_WL0_XI2.XI43.MM18_d N_XI2.XI43.NET031_XI2.XI43.MM18_g
+ N_VDD_XI2.XI43.MM18_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI53.MM18 N_WL2_XI2.XI53.MM18_d N_XI2.XI53.NET031_XI2.XI53.MM18_g
+ N_VDD_XI2.XI53.MM18_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI55.MM18 N_WL4_XI2.XI55.MM18_d N_XI2.XI55.NET031_XI2.XI55.MM18_g
+ N_VDD_XI2.XI55.MM18_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI57.MM18 N_WL6_XI2.XI57.MM18_d N_XI2.XI57.NET031_XI2.XI57.MM18_g
+ N_VDD_XI2.XI57.MM18_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI43.MM18@4 N_WL0_XI2.XI43.MM18@4_d N_XI2.XI43.NET031_XI2.XI43.MM18@4_g
+ N_VDD_XI2.XI43.MM18@4_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI53.MM18@4 N_WL2_XI2.XI53.MM18@4_d N_XI2.XI53.NET031_XI2.XI53.MM18@4_g
+ N_VDD_XI2.XI53.MM18@4_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI55.MM18@4 N_WL4_XI2.XI55.MM18@4_d N_XI2.XI55.NET031_XI2.XI55.MM18@4_g
+ N_VDD_XI2.XI55.MM18@4_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI57.MM18@4 N_WL6_XI2.XI57.MM18@4_d N_XI2.XI57.NET031_XI2.XI57.MM18@4_g
+ N_VDD_XI2.XI57.MM18@4_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI43.MM18@3 N_WL0_XI2.XI43.MM18@3_d N_XI2.XI43.NET031_XI2.XI43.MM18@3_g
+ N_VDD_XI2.XI43.MM18@3_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI53.MM18@3 N_WL2_XI2.XI53.MM18@3_d N_XI2.XI53.NET031_XI2.XI53.MM18@3_g
+ N_VDD_XI2.XI53.MM18@3_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI55.MM18@3 N_WL4_XI2.XI55.MM18@3_d N_XI2.XI55.NET031_XI2.XI55.MM18@3_g
+ N_VDD_XI2.XI55.MM18@3_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI57.MM18@3 N_WL6_XI2.XI57.MM18@3_d N_XI2.XI57.NET031_XI2.XI57.MM18@3_g
+ N_VDD_XI2.XI57.MM18@3_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI43.MM18@2 N_WL0_XI2.XI43.MM18@2_d N_XI2.XI43.NET031_XI2.XI43.MM18@2_g
+ N_VDD_XI2.XI43.MM18@2_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI53.MM18@2 N_WL2_XI2.XI53.MM18@2_d N_XI2.XI53.NET031_XI2.XI53.MM18@2_g
+ N_VDD_XI2.XI53.MM18@2_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI55.MM18@2 N_WL4_XI2.XI55.MM18@2_d N_XI2.XI55.NET031_XI2.XI55.MM18@2_g
+ N_VDD_XI2.XI55.MM18@2_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI57.MM18@2 N_WL6_XI2.XI57.MM18@2_d N_XI2.XI57.NET031_XI2.XI57.MM18@2_g
+ N_VDD_XI2.XI57.MM18@2_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI0.XI33.MM7 N_XI0.NET36_XI0.XI33.MM7_d N_XI0.NET016_XI0.XI33.MM7_g
+ N_X240.noxref_55_XI0.XI33.MM7_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI33.MM5 N_X240.noxref_55_XI0.XI33.MM5_d N_NET47_XI0.XI33.MM5_g
+ N_VSS_XI0.XI33.MM5_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI26.MM5 N_XI0.XI26.NET4_XI0.XI26.MM5_d N_XI0.NET36_XI0.XI26.MM5_g
+ N_VSS_XI0.XI26.MM5_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI23.MM5 N_XI0.XI23.NET4_XI0.XI23.MM5_d N_NET38_XI0.XI23.MM5_g
+ N_VSS_XI0.XI23.MM5_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI33.MM4 N_X240.noxref_56_XI0.XI33.MM4_d N_NET48_XI0.XI33.MM4_g
+ N_VSS_XI0.XI33.MM4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI33.MM6 N_XI0.NET36_XI0.XI33.MM6_d N_XI0.XI33.~A_XI0.XI33.MM6_g
+ N_X240.noxref_56_XI0.XI33.MM6_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI26.MM7 N_XI0.XI26.NET8_XI0.XI26.MM7_d N_XI0.XI26.NET4_XI0.XI26.MM7_g
+ N_XI0.XI26.NET31_XI0.XI26.MM7_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI0.XI23.MM7 N_XI0.XI23.NET8_XI0.XI23.MM7_d N_XI0.XI23.NET4_XI0.XI23.MM7_g
+ N_XI0.XI23.NET31_XI0.XI23.MM7_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI0.XI26.MM6 N_XI0.XI26.NET31_XI0.XI26.MM6_d N_CLK_XI0.XI26.MM6_g
+ N_VSS_XI0.XI26.MM6_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI0.XI23.MM6 N_XI0.XI23.NET31_XI0.XI23.MM6_d N_CLK_XI0.XI23.MM6_g
+ N_VSS_XI0.XI23.MM6_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI0.XI33.XI0.MM0 N_XI0.XI33.~A_XI0.XI33.XI0.MM0_d
+ N_XI0.NET016_XI0.XI33.XI0.MM0_g N_VSS_XI0.XI33.XI0.MM0_s N_VSS_XI0.XI33.MM7_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI26.MM8 N_NET48_XI0.XI26.MM8_d N_CLK_XI0.XI26.MM8_g
+ N_XI0.XI26.NET30_XI0.XI26.MM8_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI0.XI23.MM8 N_NET38_XI0.XI23.MM8_d N_CLK_XI0.XI23.MM8_g
+ N_XI0.XI23.NET30_XI0.XI23.MM8_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI0.XI26.MM10 N_XI0.XI26.NET30_XI0.XI26.MM10_d N_XI0.XI26.NET8_XI0.XI26.MM10_g
+ N_VSS_XI0.XI26.MM10_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=1.3125e-13 PD=2.5e-07 PS=5.25e-07
mXI0.XI23.MM10 N_XI0.XI23.NET30_XI0.XI23.MM10_d N_XI0.XI23.NET8_XI0.XI23.MM10_g
+ N_VSS_XI0.XI23.MM10_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=1.3125e-13 PD=2.5e-07 PS=5.25e-07
mXI0.XI26.MM9 N_NET47_XI0.XI26.MM9_d N_NET48_XI0.XI26.MM9_g N_VSS_XI0.XI26.MM9_s
+ N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.3125e-13
+ PD=1.48e-06 PS=5.25e-07
mXI0.XI32.MM4 N_XI0.NET016_XI0.XI32.MM4_d N_NET38_XI0.XI32.MM4_g
+ N_VSS_XI0.XI32.MM4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI23.MM9 N_NET37_XI0.XI23.MM9_d N_NET38_XI0.XI23.MM9_g N_VSS_XI0.XI23.MM9_s
+ N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.3125e-13
+ PD=1.48e-06 PS=5.25e-07
mXI0.XI32.MM0 N_XI0.NET016_XI0.XI32.MM0_d N_NET39_XI0.XI32.MM0_g
+ N_VSS_XI0.XI32.MM0_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI37.MM5 N_XI0.XI37.NET014_XI0.XI37.MM5_d N_XI0.NET016_XI0.XI37.MM5_g
+ N_VSS_XI0.XI37.MM5_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI32.MM1 N_XI0.NET016_XI0.XI32.MM1_d N_NET45_XI0.XI32.MM1_g
+ N_VSS_XI0.XI32.MM1_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI34.MM3 N_XI0.XI34.NET019_XI0.XI34.MM3_d N_NET47_XI0.XI34.MM3_g
+ N_VSS_XI0.XI34.MM3_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI37.MM3 N_XI0.XI37.NET37_XI0.XI37.MM3_d N_NET47_XI0.XI37.MM3_g
+ N_XI0.XI37.NET014_XI0.XI37.MM3_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI29.MM7 N_XI0.NET9_XI0.XI29.MM7_d N_NET39_XI0.XI29.MM7_g
+ N_X240.noxref_64_XI0.XI29.MM7_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI34.MM2 N_XI0.NET038_XI0.XI34.MM2_d N_XI0.NET016_XI0.XI34.MM2_g
+ N_XI0.XI34.NET019_XI0.XI34.MM2_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.397e-13 AS=1.1985e-13 PD=1.49e-06 PS=5.1e-07
mXI0.XI37.MM2 N_XI0.NET045_XI0.XI37.MM2_d N_NET46_XI0.XI37.MM2_g
+ N_XI0.XI37.NET37_XI0.XI37.MM2_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI29.MM5 N_X240.noxref_64_XI0.XI29.MM5_d N_NET38_XI0.XI29.MM5_g
+ N_VSS_XI0.XI29.MM5_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI25.MM9 N_NET43_XI0.XI25.MM9_d N_NET45_XI0.XI25.MM9_g N_VSS_XI0.XI25.MM9_s
+ N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.3125e-13
+ PD=1.48e-06 PS=5.25e-07
mXI0.XI29.MM4 N_X240.noxref_65_XI0.XI29.MM4_d N_NET37_XI0.XI29.MM4_g
+ N_VSS_XI0.XI29.MM4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI25.MM10 N_XI0.XI25.NET30_XI0.XI25.MM10_d N_XI0.XI25.NET8_XI0.XI25.MM10_g
+ N_VSS_XI0.XI25.MM10_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=1.3125e-13 PD=2.5e-07 PS=5.25e-07
mXI0.XI29.MM6 N_XI0.NET9_XI0.XI29.MM6_d N_NET41_XI0.XI29.MM6_g
+ N_X240.noxref_65_XI0.XI29.MM6_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI25.MM8 N_NET45_XI0.XI25.MM8_d N_CLK_XI0.XI25.MM8_g
+ N_XI0.XI25.NET30_XI0.XI25.MM8_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI0.XI35.XI0.MM0 N_XI0.XI35.~A_XI0.XI35.XI0.MM0_d
+ N_XI0.NET038_XI0.XI35.XI0.MM0_g N_VSS_XI0.XI35.XI0.MM0_s N_VSS_XI0.XI33.MM7_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI38.XI0.MM0 N_XI0.XI38.~A_XI0.XI38.XI0.MM0_d
+ N_XI0.NET045_XI0.XI38.XI0.MM0_g N_VSS_XI0.XI38.XI0.MM0_s N_VSS_XI0.XI33.MM7_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI25.MM6 N_XI0.XI25.NET31_XI0.XI25.MM6_d N_CLK_XI0.XI25.MM6_g
+ N_VSS_XI0.XI25.MM6_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI0.XI35.MM6 N_XI0.NET041_XI0.XI35.MM6_d N_XI0.XI35.~A_XI0.XI35.MM6_g
+ N_X240.noxref_68_XI0.XI35.MM6_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI38.MM6 N_XI0.NET049_XI0.XI38.MM6_d N_XI0.XI38.~A_XI0.XI38.MM6_g
+ N_X240.noxref_69_XI0.XI38.MM6_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI25.MM7 N_XI0.XI25.NET8_XI0.XI25.MM7_d N_XI0.XI25.NET4_XI0.XI25.MM7_g
+ N_XI0.XI25.NET31_XI0.XI25.MM7_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI0.XI35.MM4 N_X240.noxref_68_XI0.XI35.MM4_d N_NET46_XI0.XI35.MM4_g
+ N_VSS_XI0.XI35.MM4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI38.MM4 N_X240.noxref_69_XI0.XI38.MM4_d N_NET42_XI0.XI38.MM4_g
+ N_VSS_XI0.XI38.MM4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI24.MM5 N_XI0.XI24.NET4_XI0.XI24.MM5_d N_XI0.NET9_XI0.XI24.MM5_g
+ N_VSS_XI0.XI24.MM5_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI35.MM5 N_X240.noxref_70_XI0.XI35.MM5_d N_NET44_XI0.XI35.MM5_g
+ N_VSS_XI0.XI35.MM5_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI38.MM5 N_X240.noxref_71_XI0.XI38.MM5_d N_NET40_XI0.XI38.MM5_g
+ N_VSS_XI0.XI38.MM5_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI25.MM5 N_XI0.XI25.NET4_XI0.XI25.MM5_d N_XI0.NET16_XI0.XI25.MM5_g
+ N_VSS_XI0.XI25.MM5_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI35.MM7 N_XI0.NET041_XI0.XI35.MM7_d N_XI0.NET038_XI0.XI35.MM7_g
+ N_X240.noxref_70_XI0.XI35.MM7_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI38.MM7 N_XI0.NET049_XI0.XI38.MM7_d N_XI0.NET045_XI0.XI38.MM7_g
+ N_X240.noxref_71_XI0.XI38.MM7_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI24.MM7 N_XI0.XI24.NET8_XI0.XI24.MM7_d N_XI0.XI24.NET4_XI0.XI24.MM7_g
+ N_XI0.XI24.NET31_XI0.XI24.MM7_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI0.XI24.MM6 N_XI0.XI24.NET31_XI0.XI24.MM6_d N_CLK_XI0.XI24.MM6_g
+ N_VSS_XI0.XI24.MM6_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI0.XI24.MM8 N_NET39_XI0.XI24.MM8_d N_CLK_XI0.XI24.MM8_g
+ N_XI0.XI24.NET30_XI0.XI24.MM8_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI0.XI31.MM7 N_XI0.NET16_XI0.XI31.MM7_d N_XI0.NET14_XI0.XI31.MM7_g
+ N_X240.noxref_74_XI0.XI31.MM7_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI24.MM10 N_XI0.XI24.NET30_XI0.XI24.MM10_d N_XI0.XI24.NET8_XI0.XI24.MM10_g
+ N_VSS_XI0.XI24.MM10_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=1.3125e-13 PD=2.5e-07 PS=5.25e-07
mXI0.XI36.MM5 N_XI0.XI36.NET4_XI0.XI36.MM5_d N_XI0.NET041_XI0.XI36.MM5_g
+ N_VSS_XI0.XI36.MM5_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI27.MM5 N_XI0.XI27.NET4_XI0.XI27.MM5_d N_XI0.NET049_XI0.XI27.MM5_g
+ N_VSS_XI0.XI27.MM5_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI31.MM5 N_X240.noxref_74_XI0.XI31.MM5_d N_NET45_XI0.XI31.MM5_g
+ N_VSS_XI0.XI31.MM5_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI24.MM9 N_NET41_XI0.XI24.MM9_d N_NET39_XI0.XI24.MM9_g N_VSS_XI0.XI24.MM9_s
+ N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.3125e-13
+ PD=1.48e-06 PS=5.25e-07
mXI0.XI31.MM4 N_X240.noxref_75_XI0.XI31.MM4_d N_NET43_XI0.XI31.MM4_g
+ N_VSS_XI0.XI31.MM4_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI36.MM7 N_XI0.XI36.NET8_XI0.XI36.MM7_d N_XI0.XI36.NET4_XI0.XI36.MM7_g
+ N_XI0.XI36.NET31_XI0.XI36.MM7_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI0.XI27.MM7 N_XI0.XI27.NET8_XI0.XI27.MM7_d N_XI0.XI27.NET4_XI0.XI27.MM7_g
+ N_XI0.XI27.NET31_XI0.XI27.MM7_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI0.XI31.MM6 N_XI0.NET16_XI0.XI31.MM6_d N_XI0.XI31.~A_XI0.XI31.MM6_g
+ N_X240.noxref_75_XI0.XI31.MM6_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI36.MM6 N_XI0.XI36.NET31_XI0.XI36.MM6_d N_CLK_XI0.XI36.MM6_g
+ N_VSS_XI0.XI36.MM6_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI0.XI27.MM6 N_XI0.XI27.NET31_XI0.XI27.MM6_d N_CLK_XI0.XI27.MM6_g
+ N_VSS_XI0.XI27.MM6_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI0.XI30.MM3 N_XI0.XI30.NET019_XI0.XI30.MM3_d N_NET37_XI0.XI30.MM3_g
+ N_VSS_XI0.XI30.MM3_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI30.MM2 N_XI0.NET14_XI0.XI30.MM2_d N_NET41_XI0.XI30.MM2_g
+ N_XI0.XI30.NET019_XI0.XI30.MM2_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.397e-13 AS=1.1985e-13 PD=1.49e-06 PS=5.1e-07
mXI0.XI31.XI0.MM0 N_XI0.XI31.~A_XI0.XI31.XI0.MM0_d
+ N_XI0.NET14_XI0.XI31.XI0.MM0_g N_VSS_XI0.XI31.XI0.MM0_s N_VSS_XI0.XI33.MM7_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI36.MM8 N_NET44_XI0.XI36.MM8_d N_CLK_XI0.XI36.MM8_g
+ N_XI0.XI36.NET30_XI0.XI36.MM8_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI0.XI27.MM8 N_NET40_XI0.XI27.MM8_d N_CLK_XI0.XI27.MM8_g
+ N_XI0.XI27.NET30_XI0.XI27.MM8_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI0.XI36.MM10 N_XI0.XI36.NET30_XI0.XI36.MM10_d N_XI0.XI36.NET8_XI0.XI36.MM10_g
+ N_VSS_XI0.XI36.MM10_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=1.3125e-13 PD=2.5e-07 PS=5.25e-07
mXI0.XI27.MM10 N_XI0.XI27.NET30_XI0.XI27.MM10_d N_XI0.XI27.NET8_XI0.XI27.MM10_g
+ N_VSS_XI0.XI27.MM10_s N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=1.3125e-13 PD=2.5e-07 PS=5.25e-07
mXI0.XI36.MM9 N_NET46_XI0.XI36.MM9_d N_NET44_XI0.XI36.MM9_g N_VSS_XI0.XI36.MM9_s
+ N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.3125e-13
+ PD=1.48e-06 PS=5.25e-07
mXI0.XI27.MM9 N_NET42_XI0.XI27.MM9_d N_NET40_XI0.XI27.MM9_g N_VSS_XI0.XI27.MM9_s
+ N_VSS_XI0.XI33.MM7_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.3125e-13
+ PD=1.48e-06 PS=5.25e-07
mXI0.XI33.MM2 N_XI0.NET36_XI0.XI33.MM2_d N_XI0.NET016_XI0.XI33.MM2_g
+ N_X240.noxref_19_XI0.XI33.MM2_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI26.MM0 N_XI0.XI26.NET32_XI0.XI26.MM0_d N_XI0.NET36_XI0.XI26.MM0_g
+ N_VDD_XI0.XI26.MM0_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07 AD=1.125e-13
+ AS=4.5e-13 PD=2.5e-07 PS=1.9e-06
mXI0.XI23.MM0 N_XI0.XI23.NET32_XI0.XI23.MM0_d N_NET38_XI0.XI23.MM0_g
+ N_VDD_XI0.XI23.MM0_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=9e-07 AD=1.125e-13
+ AS=4.5e-13 PD=2.5e-07 PS=1.9e-06
mXI0.XI26.MM1 N_XI0.XI26.NET4_XI0.XI26.MM1_d N_CLK_XI0.XI26.MM1_g
+ N_XI0.XI26.NET32_XI0.XI26.MM1_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07
+ AD=4.41e-13 AS=1.125e-13 PD=1.88e-06 PS=2.5e-07
mXI0.XI33.MM3 N_XI0.NET36_XI0.XI33.MM3_d N_NET47_XI0.XI33.MM3_g
+ N_X240.noxref_19_XI0.XI33.MM3_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI23.MM1 N_XI0.XI23.NET4_XI0.XI23.MM1_d N_CLK_XI0.XI23.MM1_g
+ N_XI0.XI23.NET32_XI0.XI23.MM1_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=9e-07
+ AD=4.41e-13 AS=1.125e-13 PD=1.88e-06 PS=2.5e-07
mXI0.XI33.MM1 N_X240.noxref_19_XI0.XI33.MM1_d N_NET48_XI0.XI33.MM1_g
+ N_VDD_XI0.XI33.MM1_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI26.MM2 N_XI0.XI26.NET8_XI0.XI26.MM2_d N_CLK_XI0.XI26.MM2_g
+ N_VDD_XI0.XI26.MM2_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07 AD=4.59e-13
+ AS=4.41e-13 PD=1.92e-06 PS=1.88e-06
mXI0.XI33.MM0 N_X240.noxref_19_XI0.XI33.MM0_d N_XI0.XI33.~A_XI0.XI33.MM0_g
+ N_VDD_XI0.XI33.MM0_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI23.MM2 N_XI0.XI23.NET8_XI0.XI23.MM2_d N_CLK_XI0.XI23.MM2_g
+ N_VDD_XI0.XI23.MM2_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=9e-07 AD=4.59e-13
+ AS=4.41e-13 PD=1.92e-06 PS=1.88e-06
mXI0.XI26.MM3 N_NET48_XI0.XI26.MM3_d N_XI0.XI26.NET8_XI0.XI26.MM3_g
+ N_VDD_XI0.XI26.MM3_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07 AD=4.41e-13
+ AS=2.295e-13 PD=1.88e-06 PS=5.1e-07
mXI0.XI33.XI0.MM1 N_XI0.XI33.~A_XI0.XI33.XI0.MM1_d
+ N_XI0.NET016_XI0.XI33.XI0.MM1_g N_VDD_XI0.XI33.XI0.MM1_s N_VDD_XI0.XI33.MM2_b
+ P_18 L=1.8e-07 W=9.5e-07 AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI23.MM3 N_NET38_XI0.XI23.MM3_d N_XI0.XI23.NET8_XI0.XI23.MM3_g
+ N_VDD_XI0.XI23.MM3_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=9e-07 AD=4.41e-13
+ AS=2.295e-13 PD=1.88e-06 PS=5.1e-07
mXI0.XI26.MM11 N_NET48_XI0.XI26.MM11_d N_RST_XI0.XI26.MM11_g
+ N_VDD_XI0.XI26.MM11_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07 AD=2.34e-13
+ AS=2.295e-13 PD=5.2e-07 PS=5.1e-07
mXI0.XI23.MM11 N_NET38_XI0.XI23.MM11_d N_RST_XI0.XI23.MM11_g
+ N_VDD_XI0.XI23.MM11_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=9e-07 AD=2.34e-13
+ AS=2.295e-13 PD=5.2e-07 PS=5.1e-07
mXI0.XI26.MM11@2 N_NET48_XI0.XI26.MM11@2_d N_RST_XI0.XI26.MM11@2_g
+ N_VDD_XI0.XI26.MM11@2_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07
+ AD=2.34e-13 AS=2.295e-13 PD=5.2e-07 PS=5.1e-07
mXI0.XI23.MM11@2 N_NET38_XI0.XI23.MM11@2_d N_RST_XI0.XI23.MM11@2_g
+ N_VDD_XI0.XI23.MM11@2_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=9e-07
+ AD=2.34e-13 AS=2.295e-13 PD=5.2e-07 PS=5.1e-07
mXI0.XI26.MM4 N_NET47_XI0.XI26.MM4_d N_NET48_XI0.XI26.MM4_g N_VDD_XI0.XI26.MM4_s
+ N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07 AD=4.41e-13 AS=2.295e-13
+ PD=1.88e-06 PS=5.1e-07
mXI0.XI32.MM2 N_XI0.NET016_XI0.XI32.MM2_d N_NET38_XI0.XI32.MM2_g
+ N_XI0.XI32.NET36_XI0.XI32.MM2_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=2.4225e-13 PD=1.93e-06 PS=5.1e-07
mXI0.XI23.MM4 N_NET37_XI0.XI23.MM4_d N_NET38_XI0.XI23.MM4_g N_VDD_XI0.XI23.MM4_s
+ N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=9e-07 AD=4.41e-13 AS=2.295e-13
+ PD=1.88e-06 PS=5.1e-07
mXI0.XI32.MM3 N_XI0.XI32.NET36_XI0.XI32.MM3_d N_NET39_XI0.XI32.MM3_g
+ N_XI0.XI32.NET37_XI0.XI32.MM3_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9.5e-07
+ AD=2.4225e-13 AS=2.4225e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI37.MM4 N_XI0.NET045_XI0.XI37.MM4_d N_XI0.NET016_XI0.XI37.MM4_g
+ N_VDD_XI0.XI37.MM4_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI32.MM5 N_XI0.XI32.NET37_XI0.XI32.MM5_d N_NET45_XI0.XI32.MM5_g
+ N_VDD_XI0.XI32.MM5_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9.5e-07
+ AD=2.4225e-13 AS=4.655e-13 PD=5.1e-07 PS=1.93e-06
mXI0.XI34.MM0 N_XI0.NET038_XI0.XI34.MM0_d N_NET47_XI0.XI34.MM0_g
+ N_VDD_XI0.XI34.MM0_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI37.MM0 N_XI0.NET045_XI0.XI37.MM0_d N_NET47_XI0.XI37.MM0_g
+ N_VDD_XI0.XI37.MM0_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI29.MM2 N_XI0.NET9_XI0.XI29.MM2_d N_NET39_XI0.XI29.MM2_g
+ N_X240.noxref_23_XI0.XI29.MM2_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI34.MM1 N_XI0.NET038_XI0.XI34.MM1_d N_XI0.NET016_XI0.XI34.MM1_g
+ N_VDD_XI0.XI34.MM1_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.397e-13 PD=5.1e-07 PS=1.49e-06
mXI0.XI37.MM1 N_XI0.NET045_XI0.XI37.MM1_d N_NET46_XI0.XI37.MM1_g
+ N_VDD_XI0.XI37.MM1_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI29.MM3 N_XI0.NET9_XI0.XI29.MM3_d N_NET38_XI0.XI29.MM3_g
+ N_X240.noxref_23_XI0.XI29.MM3_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI25.MM4 N_NET43_XI0.XI25.MM4_d N_NET45_XI0.XI25.MM4_g N_VDD_XI0.XI25.MM4_s
+ N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07 AD=4.41e-13 AS=2.295e-13
+ PD=1.88e-06 PS=5.1e-07
mXI0.XI29.MM1 N_X240.noxref_23_XI0.XI29.MM1_d N_NET37_XI0.XI29.MM1_g
+ N_VDD_XI0.XI29.MM1_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI25.MM11 N_NET45_XI0.XI25.MM11_d N_RST_XI0.XI25.MM11_g
+ N_VDD_XI0.XI25.MM11_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07 AD=2.34e-13
+ AS=2.295e-13 PD=5.2e-07 PS=5.1e-07
mXI0.XI29.MM0 N_X240.noxref_23_XI0.XI29.MM0_d N_NET41_XI0.XI29.MM0_g
+ N_VDD_XI0.XI29.MM0_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI35.XI0.MM1 N_XI0.XI35.~A_XI0.XI35.XI0.MM1_d
+ N_XI0.NET038_XI0.XI35.XI0.MM1_g N_VDD_XI0.XI35.XI0.MM1_s N_VDD_XI0.XI33.MM2_b
+ P_18 L=1.8e-07 W=9.5e-07 AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI38.XI0.MM1 N_XI0.XI38.~A_XI0.XI38.XI0.MM1_d
+ N_XI0.NET045_XI0.XI38.XI0.MM1_g N_VDD_XI0.XI38.XI0.MM1_s N_VDD_XI0.XI37.MM4_b
+ P_18 L=1.8e-07 W=9.5e-07 AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI25.MM11@2 N_NET45_XI0.XI25.MM11@2_d N_RST_XI0.XI25.MM11@2_g
+ N_VDD_XI0.XI25.MM11@2_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07
+ AD=2.34e-13 AS=2.295e-13 PD=5.2e-07 PS=5.1e-07
mXI0.XI25.MM3 N_NET45_XI0.XI25.MM3_d N_XI0.XI25.NET8_XI0.XI25.MM3_g
+ N_VDD_XI0.XI25.MM3_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07 AD=4.41e-13
+ AS=2.295e-13 PD=1.88e-06 PS=5.1e-07
mXI0.XI35.MM0 N_X240.noxref_25_XI0.XI35.MM0_d N_XI0.XI35.~A_XI0.XI35.MM0_g
+ N_VDD_XI0.XI35.MM0_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI38.MM0 N_X240.noxref_26_XI0.XI38.MM0_d N_XI0.XI38.~A_XI0.XI38.MM0_g
+ N_VDD_XI0.XI38.MM0_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI24.MM0 N_XI0.XI24.NET32_XI0.XI24.MM0_d N_XI0.NET9_XI0.XI24.MM0_g
+ N_VDD_XI0.XI24.MM0_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=9e-07 AD=1.125e-13
+ AS=4.5e-13 PD=2.5e-07 PS=1.9e-06
mXI0.XI24.MM1 N_XI0.XI24.NET4_XI0.XI24.MM1_d N_CLK_XI0.XI24.MM1_g
+ N_XI0.XI24.NET32_XI0.XI24.MM1_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=9e-07
+ AD=4.41e-13 AS=1.125e-13 PD=1.88e-06 PS=2.5e-07
mXI0.XI35.MM1 N_X240.noxref_25_XI0.XI35.MM1_d N_NET46_XI0.XI35.MM1_g
+ N_VDD_XI0.XI35.MM1_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI25.MM2 N_XI0.XI25.NET8_XI0.XI25.MM2_d N_CLK_XI0.XI25.MM2_g
+ N_VDD_XI0.XI25.MM2_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07 AD=4.59e-13
+ AS=4.41e-13 PD=1.92e-06 PS=1.88e-06
mXI0.XI38.MM1 N_X240.noxref_26_XI0.XI38.MM1_d N_NET42_XI0.XI38.MM1_g
+ N_VDD_XI0.XI38.MM1_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI35.MM3 N_XI0.NET041_XI0.XI35.MM3_d N_NET44_XI0.XI35.MM3_g
+ N_X240.noxref_25_XI0.XI35.MM3_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI38.MM3 N_XI0.NET049_XI0.XI38.MM3_d N_NET40_XI0.XI38.MM3_g
+ N_X240.noxref_26_XI0.XI38.MM3_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI35.MM2 N_XI0.NET041_XI0.XI35.MM2_d N_XI0.NET038_XI0.XI35.MM2_g
+ N_X240.noxref_25_XI0.XI35.MM2_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI24.MM2 N_XI0.XI24.NET8_XI0.XI24.MM2_d N_CLK_XI0.XI24.MM2_g
+ N_VDD_XI0.XI24.MM2_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=9e-07 AD=4.59e-13
+ AS=4.41e-13 PD=1.92e-06 PS=1.88e-06
mXI0.XI38.MM2 N_XI0.NET049_XI0.XI38.MM2_d N_XI0.NET045_XI0.XI38.MM2_g
+ N_X240.noxref_26_XI0.XI38.MM2_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI25.MM1 N_XI0.XI25.NET4_XI0.XI25.MM1_d N_CLK_XI0.XI25.MM1_g
+ N_XI0.XI25.NET32_XI0.XI25.MM1_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07
+ AD=4.41e-13 AS=1.125e-13 PD=1.88e-06 PS=2.5e-07
mXI0.XI25.MM0 N_XI0.XI25.NET32_XI0.XI25.MM0_d N_XI0.NET16_XI0.XI25.MM0_g
+ N_VDD_XI0.XI25.MM0_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07 AD=1.125e-13
+ AS=4.5e-13 PD=2.5e-07 PS=1.9e-06
mXI0.XI24.MM3 N_NET39_XI0.XI24.MM3_d N_XI0.XI24.NET8_XI0.XI24.MM3_g
+ N_VDD_XI0.XI24.MM3_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=9e-07 AD=4.41e-13
+ AS=2.295e-13 PD=1.88e-06 PS=5.1e-07
mXI0.XI36.MM0 N_XI0.XI36.NET32_XI0.XI36.MM0_d N_XI0.NET041_XI0.XI36.MM0_g
+ N_VDD_XI0.XI36.MM0_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07 AD=1.125e-13
+ AS=4.5e-13 PD=2.5e-07 PS=1.9e-06
mXI0.XI24.MM11 N_NET39_XI0.XI24.MM11_d N_RST_XI0.XI24.MM11_g
+ N_VDD_XI0.XI24.MM11_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=9e-07 AD=2.34e-13
+ AS=2.295e-13 PD=5.2e-07 PS=5.1e-07
mXI0.XI27.MM0 N_XI0.XI27.NET32_XI0.XI27.MM0_d N_XI0.NET049_XI0.XI27.MM0_g
+ N_VDD_XI0.XI27.MM0_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=9e-07 AD=1.125e-13
+ AS=4.5e-13 PD=2.5e-07 PS=1.9e-06
mXI0.XI36.MM1 N_XI0.XI36.NET4_XI0.XI36.MM1_d N_CLK_XI0.XI36.MM1_g
+ N_XI0.XI36.NET32_XI0.XI36.MM1_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07
+ AD=4.41e-13 AS=1.125e-13 PD=1.88e-06 PS=2.5e-07
mXI0.XI27.MM1 N_XI0.XI27.NET4_XI0.XI27.MM1_d N_CLK_XI0.XI27.MM1_g
+ N_XI0.XI27.NET32_XI0.XI27.MM1_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=9e-07
+ AD=4.41e-13 AS=1.125e-13 PD=1.88e-06 PS=2.5e-07
mXI0.XI31.MM2 N_XI0.NET16_XI0.XI31.MM2_d N_XI0.NET14_XI0.XI31.MM2_g
+ N_X240.noxref_29_XI0.XI31.MM2_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI24.MM11@2 N_NET39_XI0.XI24.MM11@2_d N_RST_XI0.XI24.MM11@2_g
+ N_VDD_XI0.XI24.MM11@2_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=9e-07
+ AD=2.34e-13 AS=2.295e-13 PD=5.2e-07 PS=5.1e-07
mXI0.XI31.MM3 N_XI0.NET16_XI0.XI31.MM3_d N_NET45_XI0.XI31.MM3_g
+ N_X240.noxref_29_XI0.XI31.MM3_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI24.MM4 N_NET41_XI0.XI24.MM4_d N_NET39_XI0.XI24.MM4_g N_VDD_XI0.XI24.MM4_s
+ N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=9e-07 AD=4.41e-13 AS=2.295e-13
+ PD=1.88e-06 PS=5.1e-07
mXI0.XI36.MM2 N_XI0.XI36.NET8_XI0.XI36.MM2_d N_CLK_XI0.XI36.MM2_g
+ N_VDD_XI0.XI36.MM2_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07 AD=4.59e-13
+ AS=4.41e-13 PD=1.92e-06 PS=1.88e-06
mXI0.XI31.MM1 N_X240.noxref_29_XI0.XI31.MM1_d N_NET43_XI0.XI31.MM1_g
+ N_VDD_XI0.XI31.MM1_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI27.MM2 N_XI0.XI27.NET8_XI0.XI27.MM2_d N_CLK_XI0.XI27.MM2_g
+ N_VDD_XI0.XI27.MM2_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=9e-07 AD=4.59e-13
+ AS=4.41e-13 PD=1.92e-06 PS=1.88e-06
mXI0.XI31.MM0 N_X240.noxref_29_XI0.XI31.MM0_d N_XI0.XI31.~A_XI0.XI31.MM0_g
+ N_VDD_XI0.XI31.MM0_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI36.MM3 N_NET44_XI0.XI36.MM3_d N_XI0.XI36.NET8_XI0.XI36.MM3_g
+ N_VDD_XI0.XI36.MM3_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07 AD=4.41e-13
+ AS=2.295e-13 PD=1.88e-06 PS=5.1e-07
mXI0.XI27.MM3 N_NET40_XI0.XI27.MM3_d N_XI0.XI27.NET8_XI0.XI27.MM3_g
+ N_VDD_XI0.XI27.MM3_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=9e-07 AD=4.41e-13
+ AS=2.295e-13 PD=1.88e-06 PS=5.1e-07
mXI0.XI30.MM0 N_XI0.NET14_XI0.XI30.MM0_d N_NET37_XI0.XI30.MM0_g
+ N_VDD_XI0.XI30.MM0_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI36.MM11 N_NET44_XI0.XI36.MM11_d N_RST_XI0.XI36.MM11_g
+ N_VDD_XI0.XI36.MM11_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07 AD=2.34e-13
+ AS=2.295e-13 PD=5.2e-07 PS=5.1e-07
mXI0.XI27.MM11 N_NET40_XI0.XI27.MM11_d N_RST_XI0.XI27.MM11_g
+ N_VDD_XI0.XI27.MM11_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=9e-07 AD=2.34e-13
+ AS=2.295e-13 PD=5.2e-07 PS=5.1e-07
mXI0.XI30.MM1 N_XI0.NET14_XI0.XI30.MM1_d N_NET41_XI0.XI30.MM1_g
+ N_VDD_XI0.XI30.MM1_s N_VDD_XI0.XI23.MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.397e-13 PD=5.1e-07 PS=1.49e-06
mXI0.XI31.XI0.MM1 N_XI0.XI31.~A_XI0.XI31.XI0.MM1_d
+ N_XI0.NET14_XI0.XI31.XI0.MM1_g N_VDD_XI0.XI31.XI0.MM1_s N_VDD_XI0.XI33.MM2_b
+ P_18 L=1.8e-07 W=9.5e-07 AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI36.MM11@2 N_NET44_XI0.XI36.MM11@2_d N_RST_XI0.XI36.MM11@2_g
+ N_VDD_XI0.XI36.MM11@2_s N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07
+ AD=2.34e-13 AS=2.295e-13 PD=5.2e-07 PS=5.1e-07
mXI0.XI27.MM11@2 N_NET40_XI0.XI27.MM11@2_d N_RST_XI0.XI27.MM11@2_g
+ N_VDD_XI0.XI27.MM11@2_s N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=9e-07
+ AD=2.34e-13 AS=2.295e-13 PD=5.2e-07 PS=5.1e-07
mXI0.XI36.MM4 N_NET46_XI0.XI36.MM4_d N_NET44_XI0.XI36.MM4_g N_VDD_XI0.XI36.MM4_s
+ N_VDD_XI0.XI33.MM2_b P_18 L=1.8e-07 W=9e-07 AD=4.41e-13 AS=2.295e-13
+ PD=1.88e-06 PS=5.1e-07
mXI0.XI27.MM4 N_NET42_XI0.XI27.MM4_d N_NET40_XI0.XI27.MM4_g N_VDD_XI0.XI27.MM4_s
+ N_VDD_XI0.XI37.MM4_b P_18 L=1.8e-07 W=9e-07 AD=4.41e-13 AS=2.295e-13
+ PD=1.88e-06 PS=5.1e-07
*
.include "/home/IC/final/READ/read_out.pex.spi.READ_OUT.pxi"
*
.ends
*
*
